------------------------------------------------------------------------
-- Script created table file
------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library DSO;
use DSO.Global.all;

package pFirCoeff is
constant cFirCoeff : aInputValues(0 to 128-1) := ( 473, -176, -5998, 25855, 44407, 4289, -4569, 1254, 1254, -4569, 4289, 44407, 25855, -5998, -176, 473, 223, 314, -3444, 10120, 23194, 4584, -3041, 764, 520, -634, -2493, 15827, 20534, 197, -1899, 770, 770, -1899, 197, 20534, 15827, -2493, -634, 520, 764, -3041, 4584, 23194, 10120, -3444, 314, 223, -446, 88, 7313, 6625, -299, 0, 0, 0, -577, 576, 7898, 5860, -587, 0, 0, 0, -703, 1161, 8358, 5044, -779, 0, 0, 0, -811, 1832, 8674, 4207, -885, 0, 0, 0, -887, 2577, 8836, 3376, -916, 0, 0, 0, -916, 3376, 8836, 2577, -887, 0, 0, 0, -885, 4207, 8674, 1832, -811, 0, 0, 0, -779, 5044, 8358, 1161, -703, 0, 0, 0, -587, 5860, 7898, 576, -577, 0, 0, 0, -299, 6625, 7313, 88, -446, 0, 0, 0);
end;
