------------------------------------------------------------------------
-- Script created table file
------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library DSO;
use DSO.Global.all;

package pLongInputValues is
constant cLongInputValues : aInputValues(0 to 6000-1) := ( 10127, 11528, 2440, 12226, 9140, 2994, 5479, 9018, 14272, 14663, 5231, 15337, 15477, 10090, 14189, 6552, 10228, 16485, 15297, 17615, 14253, 7077, 17185, 18508, 15729, 16981, 17104, 13171, 16644, 11102, 17849, 10016, 13268, 10782, 11693, 20746, 19491, 15231, 23159, 12410, 17579, 17182, 22104, 22754, 15710, 19653, 19410, 22120, 23170, 24005, 18521, 23676, 23666, 18013, 17773, 22632, 28480, 21295, 24531, 20454, 27096, 21394, 24698, 27306, 29898, 31000, 26308, 21658, 22062, 23641, 30948, 24149, 31174, 24563, 33102, 26387, 24806, 25731, 30398, 28943, 27742, 33784, 31086, 30920, 35612, 28259, 34202, 34419, 30175, 32691, 27014, 27004, 33008, 36255, 38373, 28927, 34469, 33518, 28248, 32415, 30550, 38416, 32833, 35695, 31559, 37060, 33209, 38162, 38821, 39766, 36410, 32220, 34200, 42682, 33734, 42081, 38840, 44584, 33738, 38355, 34524, 45055, 33730, 43234, 43960, 44794, 35549, 39563, 38085, 44807, 40569, 46553, 37969, 39159, 37935, 38020, 47060, 43764, 43600, 38912, 47642, 45048, 41968, 44113, 42956, 39212, 41372, 40148, 41059, 41914, 44230, 39973, 50433, 51113, 45811, 45961, 44302, 51249, 45013, 42065, 50294, 45745, 44118, 46231, 42679, 43260, 53180, 53500, 49055, 42987, 45242, 46813, 52599, 43023, 43494, 45150, 51074, 52204, 51323, 49079, 50366, 47470, 53001, 46423, 52547, 46598, 48946, 52162, 54141, 45823, 56163, 54418, 51042, 50533, 50768, 49177, 51714, 51840, 55636, 55456, 53734, 50621, 55931, 52657, 50546, 57723, 57045, 53196, 54147, 53796, 49296, 50496, 52613, 49783, 57251, 49484, 49923, 49319, 50065, 52632, 51185, 58622, 52727, 49819, 58550, 59499, 53021, 49112, 50925, 52780, 55062, 51086, 55227, 56565, 50692, 49462, 51649, 51939, 53232, 54261, 49186, 51336, 57844, 48550, 59409, 57023, 54115, 55204, 51093, 53765, 59844, 54822, 54508, 51010, 54104, 55723, 56375, 52941, 52586, 60050, 48572, 58769, 59084, 57646, 49209, 51146, 52001, 56120, 49536, 56549, 49100, 55655, 53688, 57079, 56260, 58487, 58283, 51517, 55859, 49763, 47689, 56233, 53229, 52923, 57980, 54357, 54383, 57227, 56504, 53671, 48846, 49456, 57172, 46747, 52224, 48257, 57945, 54649, 51999, 51552, 46496, 53904, 46094, 46344, 51671, 46444, 55037, 54923, 53667, 46652, 52686, 50872, 56235, 52210, 53916, 49616, 49235, 53848, 44777, 45248, 45603, 48094, 53272, 52799, 43704, 47651, 49050, 47581, 50332, 49838, 45640, 47176, 42008, 53535, 43531, 42641, 45694, 43434, 46790, 44818, 52036, 51493, 40865, 48959, 43137, 44819, 46154, 50742, 44235, 50874, 42477, 47115, 46514, 44797, 46529, 45962, 39884, 39091, 49403, 39227, 37363, 43541, 47211, 44448, 38476, 40427, 41331, 47409, 37253, 45476, 42726, 39279, 36833, 39483, 39918, 35345, 40782, 36184, 37875, 40047, 35832, 36075, 39790, 35322, 41837, 43518, 40245, 35355, 38020, 32044, 41439, 40882, 39899, 32945, 36729, 29593, 34208, 32609, 30542, 30506, 33204, 28994, 34827, 33039, 35502, 35299, 34307, 26759, 26929, 29698, 31989, 33222, 29987, 34700, 33214, 35971, 30435, 27686, 24775, 30603, 32361, 27809, 23530, 25380, 23750, 25015, 26662, 27439, 26326, 31092, 26508, 31365, 27400, 30981, 22058, 27030, 22083, 26418, 26419, 18575, 20546, 19892, 24960, 26805, 20492, 25464, 23910, 15561, 22454, 19568, 25661, 14341, 19614, 18864, 19014, 22452, 16762, 22043, 17972, 12426, 13822, 20110, 16822, 12659, 14635, 17550, 12241, 18536, 12264, 20100, 11984, 17672, 10418, 11311, 8644, 14194, 15186, 13237, 11479, 13816, 13553, 13631, 12808, 16238, 7058, 12790, 6784, 5073, 10654, 8456, 8257, 10405, 11409, 6041, 9498, 6230, 11061, 10649, 3395, 7397, 6718, 5914, 9581, 1981, 2320, -380, 9212, 5361, 3055, 4680, 3237, 4172, 2623, 4457, 1761, 7141, -2505, -4168, -4422, -5278, -1467, -1239, -2535, 1961, 26, 1464, 3105, 3288, -6424, -7363, -940, -8501, -3594, -3831, -138, -4971, -6368, -3311, -2763, -5724, -8095, -10772, -5806, -10004, -12920, -4644, -11110, -8992, -6323, -10573, -6314, -10720, -7526, -7563, -11005, -16387, -12918, -12074, -14214, -15379, -8129, -13134, -7893, -14160, -9881, -14649, -9961, -10882, -15711, -17932, -11279, -9636, -17405, -13532, -16608, -12116, -13164, -20686, -12576, -11300, -17298, -13103, -16938, -22425, -22142, -19906, -16044, -15375, -16062, -22003, -19660, -25269, -25260, -25216, -18927, -21390, -25322, -21889, -26325, -27687, -18337, -22079, -17871, -20921, -22535, -19969, -19439, -18351, -30504, -20309, -23591, -19272, -25077, -25887, -22234, -29376, -26343, -21710, -25866, -22826, -24331, -26391, -30699, -25855, -33099, -26771, -26562, -25943, -24211, -23315, -26094, -28561, -24582, -28984, -35975, -34922, -26175, -30935, -26782, -34639, -30696, -29952, -37351, -30512, -33741, -37699, -32576, -36340, -37358, -36543, -37431, -37094, -39034, -32062, -36493, -33567, -31847, -34378, -34100, -35356, -39391, -35133, -30918, -30823, -38256, -39155, -35008, -34250, -37091, -39783, -30981, -41565, -41422, -41124, -40968, -35624, -36329, -42752, -32284, -34856, -34873, -43132, -33646, -32877, -32395, -34028, -35030, -38428, -42591, -40039, -43341, -44692, -33848, -41644, -41817, -41468, -39951, -37865, -45473, -35716, -39224, -35757, -41950, -40853, -45663, -44265, -38490, -42573, -35807, -45292, -34873, -40353, -38411, -34952, -43600, -42138, -41594, -38049, -37454, -46170, -45286, -43151, -46856, -41297, -43589, -45567, -45210, -36858, -39669, -42203, -36890, -46670, -38968, -39111, -41243, -45825, -40870, -44479, -46500, -45574, -37364, -47310, -45262, -47550, -42882, -48057, -37405, -45857, -47105, -44526, -42732, -47003, -36221, -44213, -44623, -47450, -44589, -47612, -42061, -38956, -40508, -47011, -47096, -38674, -37104, -41553, -46641, -37966, -43812, -44307, -38814, -47648, -47145, -39631, -40362, -41246, -38741, -38960, -38012, -43906, -38970, -40548, -42418, -46393, -37663, -42933, -39605, -37926, -45528, -45175, -40014, -40712, -35745, -36767, -37462, -45613, -45266, -44988, -36338, -34501, -37533, -44088, -36868, -44152, -43964, -37551, -41207, -37181, -35923, -37813, -35809, -41787, -35640, -32681, -33812, -43104, -39603, -39445, -35510, -36432, -33994, -38947, -40763, -42067, -33667, -40357, -38015, -35902, -39651, -34526, -36278, -40140, -32392, -40456, -37970, -38498, -34802, -39942, -35998, -39460, -39207, -30937, -36714, -32784, -28263, -34506, -31171, -30233, -33981, -31117, -37518, -27402, -36219, -35086, -28491, -32045, -28464, -32772, -34065, -36715, -28851, -31595, -31130, -29026, -35463, -32170, -26458, -27174, -33855, -33590, -33838, -34648, -29429, -26414, -25388, -27485, -32362, -25839, -31712, -31398, -31607, -30860, -30320, -29757, -28068, -27853, -28816, -28182, -20210, -22265, -23809, -28051, -27482, -28868, -18543, -20800, -22355, -25059, -26591, -20844, -16192, -25803, -24501, -22576, -26218, -18611, -21755, -14503, -21250, -18360, -23726, -20732, -23129, -15671, -14048, -20061, -15762, -20219, -17103, -13199, -15765, -18660, -18827, -16709, -16801, -17290, -14623, -12129, -15693, -15359, -18756, -19692, -16211, -15604, -11273, -7338, -7314, -12796, -15137, -8544, -8317, -8260, -7940, -15346, -8120, -10467, -13208, -14292, -5262, -12794, -12644, -6296, -3253, -7518, -4983, -11313, -1376, -6059, -4092, -11554, -1944, -2380, -9663, -4486, -6593, -3636, -5119, -4627, -7156, -5958, -8492, 2696, -261, 3401, -5574, 3861, 2636, 316, -1040, -2939, 3323, -2686, -4368, 4412, 3554, 4387, 3807, 1420, 1381, 6813, 1102, 7398, 7394, 8459, 4582, 6453, 10557, 4747, 421, 10451, 7914, 4888, 12931, 3915, 9382, 9113, 6790, 4138, 3029, 8106, 5551, 12385, 8401, 14385, 13392, 11726, 7275, 16988, 8944, 17194, 9044, 11150, 8001, 14964, 9723, 8388, 16863, 12631, 16706, 13667, 16900, 9894, 20909, 19879, 19515, 20622, 15734, 18850, 18640, 18386, 15605, 15579, 18319, 15911, 23156, 25638, 14399, 20786, 15666, 24576, 27120, 16287, 27094, 16272, 24584, 26073, 23348, 27866, 28314, 25303, 19699, 20944, 20794, 19381, 20445, 26866, 31041, 24260, 25213, 32406, 32212, 29242, 33272, 30873, 25957, 30154, 25379, 26266, 31172, 29601, 28464, 31032, 33078, 31327, 31206, 31849, 31244, 26326, 34264, 37856, 30375, 38065, 30785, 37549, 32593, 32346, 30235, 29373, 31829, 37106, 38035, 37204, 29199, 39489, 40683, 39097, 30553, 34835, 39003, 39541, 33682, 34453, 39555, 37426, 39417, 34974, 34484, 42577, 42043, 44285, 34538, 35654, 34869, 39796, 36436, 45122, 35726, 35275, 41672, 44475, 39128, 37730, 39863, 38512, 42331, 47308, 44161, 37999, 41683, 37822, 43401, 42753, 49765, 47711, 43967, 49081, 40138, 43364, 50024, 50084, 47802, 46830, 43688, 51008, 41397, 48871, 48025, 50442, 45363, 49765, 50957, 44934, 47863, 53167, 48139, 45653, 49290, 46320, 51242, 47257, 48348, 50932, 54426, 46789, 53078, 52024, 54753, 43765, 47815, 51632, 47164, 46674, 52596, 51675, 51387, 52349, 45076, 48824, 50175, 47750, 53578, 55389, 48566, 54092, 47042, 55572, 47254, 52773, 50192, 55600, 52039, 51959, 56720, 50490, 51737, 58019, 46993, 58295, 48922, 54761, 53863, 55005, 51288, 54483, 56852, 47368, 48211, 59015, 55174, 50166, 52299, 48959, 50777, 50699, 51638, 49521, 51926, 49239, 58474, 48989, 59104, 52736, 48529, 52117, 56893, 57628, 54642, 56370, 58893, 48798, 51817, 48728, 50543, 56882, 56911, 58802, 55247, 49081, 59358, 57883, 51679, 54784, 60098, 56847, 58325, 53422, 53860, 54933, 51400, 57169, 54193, 55895, 51782, 49719, 53753, 52359, 57461, 57333, 55950, 49462, 48073, 54523, 51357, 59012, 59466, 51046, 57196, 58293, 54639, 58038, 58700, 53882, 55982, 54090, 47383, 52388, 54728, 53149, 51281, 58017, 56643, 56801, 50975, 53553, 56838, 57488, 54205, 48549, 53849, 46740, 50681, 53723, 56842, 55261, 51224, 54402, 50201, 56783, 56869, 55265, 49422, 50102, 47477, 53844, 54911, 55162, 50753, 51118, 45565, 54491, 48943, 45860, 54095, 52307, 53616, 46273, 50815, 50565, 43892, 47178, 45439, 50613, 45238, 52475, 51483, 46063, 47208, 49423, 50946, 48075, 47491, 44327, 45733, 48669, 50556, 48413, 39773, 47510, 44486, 44300, 40253, 48485, 42397, 41265, 42243, 42455, 44327, 44323, 42129, 41964, 43184, 44703, 48044, 45089, 41004, 46009, 37396, 36301, 36382, 37136, 38861, 38380, 34672, 40829, 35255, 35657, 41284, 43818, 44985, 39900, 44816, 39248, 38564, 36111, 37082, 37599, 32296, 41913, 31757, 36004, 40478, 35032, 37436, 39672, 40248, 40549, 31381, 31956, 39421, 35505, 34180, 35247, 37490, 33774, 29547, 32332, 31767, 38003, 33576, 34229, 34272, 29513, 31306, 31525, 26439, 31068, 32407, 28908, 33585, 32055, 27311, 28180, 27094, 31518, 30751, 26815, 29721, 32481, 30266, 29044, 21580, 24688, 26835, 24972, 19762, 21634, 28656, 18506, 28452, 18697, 25541, 23222, 19536, 23516, 17811, 24146, 22996, 16155, 15872, 16743, 14853, 19574, 24072, 21192, 19728, 23582, 14051, 23530, 13591, 18229, 13427, 18152, 11167, 20062, 20755, 21281, 21830, 15723, 12608, 10253, 14864, 15503, 17342, 8845, 15523, 13479, 9008, 17963, 13466, 11358, 17102, 13352, 10592, 14966, 10961, 10916, 12136, 8061, 6216, 10009, 13179, 7328, 3479, 7170, 5135, 6052, 10958, 5473, 5008, 4346, 1388, 2531, 138, 3966, 1587, 1770, 3002, -986, 3244, 5489, -394, 5833, -3042, 512, -4498, -2180, -5126, -3162, -4026, -2813, -4237, -4974, 275, 3619, 3782, -5177, -2323, -3908, -2424, -5844, -8511, -4371, -7833, -9911, 990, -5625, 482, -2214, -11613, -3795, -3776, -4802, -6214, -10535, -4143, -10998, -9565, -3584, -4290, -10052, -11358, -8141, -4791, -5091, -9205, -12613, -6621, -11856, -6569, -17355, -11617, -9678, -16436, -14819, -16892, -15551, -14840, -13372, -19674, -13871, -17496, -18171, -18423, -19768, -10364, -10884, -12563, -13922, -20850, -18891, -21225, -23751, -20213, -15855, -17013, -18264, -19778, -21865, -19539, -16661, -16906, -19408, -17592, -19075, -25625, -21279, -23422, -26747, -26322, -25961, -20489, -23635, -20708, -26226, -29444, -23382, -26670, -18865, -19580, -26009, -30678, -23113, -21345, -19954, -31210, -26693, -25325, -24293, -24121, -25179, -24472, -28949, -26661, -32490, -33410, -22505, -31097, -27568, -23350, -32920, -33039, -31452, -24527, -31268, -32885, -34547, -31789, -32256, -35389, -31918, -36253, -30136, -37604, -31012, -28588, -35458, -33077, -31796, -38101, -33036, -31453, -36706, -29455, -28012, -29686, -33960, -36867, -31393, -37704, -29180, -33406, -33807, -39122, -40271, -38438, -31316, -30835, -33535, -33375, -39494, -35465, -32780, -37827, -30918, -41890, -39242, -37080, -42650, -34762, -36931, -37387, -33889, -33666, -34630, -40433, -38932, -35432, -43294, -43410, -41591, -38630, -33337, -36606, -41517, -41866, -35229, -34590, -37972, -42698, -44803, -35857, -39005, -34712, -45496, -39268, -42963, -36502, -44260, -41305, -41973, -36825, -38702, -44431, -43168, -45457, -39039, -40314, -45214, -45540, -41637, -36484, -40830, -47143, -46941, -37931, -42242, -43116, -38251, -43420, -41433, -39308, -37416, -43994, -40150, -36264, -47130, -40993, -43105, -44390, -44956, -39006, -36171, -45936, -38779, -45848, -36251, -38550, -43113, -39443, -42223, -38476, -43930, -47341, -41091, -37233, -45862, -42972, -39138, -47683, -36726, -38909, -41357, -45855, -42042, -41774, -36000, -37650, -36319, -39702, -42987, -36539, -41991, -44935, -42906, -39137, -40855, -38416, -35484, -35829, -40926, -35698, -45866, -46579, -43466, -40075, -40601, -36068, -40346, -41583, -40173, -38050, -46362, -36825, -44682, -40548, -43135, -41694, -38076, -43919, -42510, -43387, -43329, -41642, -34867, -39700, -40406, -43011, -33381, -40043, -34662, -37313, -40077, -33926, -34921, -38659, -34329, -33188, -38721, -39739, -36447, -32636, -34915, -38696, -34250, -31471, -36292, -36184, -38804, -41553, -40072, -40998, -36382, -41708, -30636, -33765, -41343, -40837, -38532, -35399, -39189, -40456, -31629, -35960, -30651, -34627, -34457, -38955, -38775, -38100, -31858, -35935, -28516, -28143, -26677, -32216, -35268, -35009, -31074, -28166, -32973, -31408, -29065, -25516, -34431, -27550, -29012, -30551, -24910, -30627, -33002, -27315, -27218, -30577, -24637, -22054, -22062, -32142, -30656, -32953, -25693, -31460, -27660, -21688, -25514, -27447, -29156, -26123, -19679, -29482, -25068, -20178, -29752, -21699, -17996, -26146, -27709, -20818, -17872, -21229, -17498, -25772, -18761, -23434, -22313, -25233, -16984, -19072, -17448, -16391, -25034, -14123, -19331, -15966, -15861, -14530, -22404, -18514, -16312, -12261, -13167, -12173, -15679, -15409, -11858, -21477, -10950, -16439, -20644, -11813, -18669, -18526, -12680, -16642, -15524, -14311, -13977, -13941, -10965, -16025, -15487, -16332, -13294, -7627, -13800, -7411, -7699, -5830, -5496, -11655, -11174, -8309, -10405, -4007, -3977, -6740, -9994, -4667, -9764, -6785, -7358, -5207, 551, -2006, 1005, -7691, -3852, -9309, -506, -2077, 1298, 3177, 2766, -3205, -7840, -1023, -4741, -4302, -2717, -5189, 2969, 3281, 1108, -1065, 5196, 2124, 7309, 6831, 666, 3258, 1152, 4784, 7182, 6873, -304, 8401, -909, 4088, 8213, 9119, 4429, 10345, 13484, 7008, 6997, 9492, 12333, 12897, 21929, 12658, 20463, 16539, 25922, 19048, 24274, 31433, 24806, 22196, 25283, 28549, 28786, 28508, 37967, 35819, 40045, 34547, 41385, 30854, 38837, 41787, 35541, 44532, 43002, 44226, 41589, 44595, 39320, 38310, 39596, 43040, 46110, 39665, 41025, 46523, 43447, 47841, 38149, 45420, 43298, 37802, 40141, 38770, 40692, 42575, 33601, 41605, 41162, 34572, 34716, 35622, 36323, 35937, 35195, 29785, 29269, 34590, 28900, 31139, 23098, 26113, 24522, 27837, 16026, 19773, 18757, 12266, 20782, 19219, 12518, 15309, 6324, 10652, 4960, 5828, 9268, 94, 33, 843, -2258, 1959, 2911, -8393, -8754, -4425, -9630, -3661, -4901, -10062, -8627, -15299, -13643, -10471, -16661, -13172, -16732, -20533, -19579, -17457, -26600, -25023, -18579, -26400, -23972, -21667, -21106, -25758, -32804, -34106, -27469, -28414, -23934, -26767, -27954, -29761, -33015, -24574, -29635, -35706, -27547, -29497, -34822, -24521, -30940, -31772, -32738, -29885, -30354, -24673, -31118, -27931, -27145, -19179, -23638, -19045, -20010, -16925, -24044, -12630, -13174, -21740, -15641, -16218, -11399, -15047, -9633, -8129, -6924, -7486, -11183, -4115, -4080, -6366, -786, 452, 3015, 7440, 7542, 10972, 2447, 5827, 10076, 17441, 16751, 14004, 13894, 11891, 21401, 19849, 17400, 21371, 19461, 27673, 24207, 32250, 22198, 33055, 31648, 31589, 33900, 35746, 29012, 39304, 29704, 33846, 33190, 42869, 33156, 39929, 41147, 41811, 44829, 35475, 44998, 41823, 44065, 38450, 42585, 44600, 47704, 41523, 37133, 36683, 43419, 45216, 43686, 39201, 46091, 40533, 45300, 34176, 35228, 41473, 42502, 40220, 33610, 31097, 38668, 37045, 29945, 28486, 28634, 33754, 32620, 28510, 27416, 22832, 26648, 26629, 21137, 19955, 18932, 15404, 18889, 20332, 19068, 15788, 8576, 12398, 4315, 2853, 2302, 394, 4330, -3198, 4481, 1938, 3051, -3495, -2849, -1306, -6823, -11172, -4044, -16588, -14284, -7650, -16119, -17901, -21248, -12709, -23129, -21735, -15857, -21556, -21024, -22234, -21627, -30430, -25113, -31741, -22758, -29189, -23589, -31293, -27662, -23731, -34776, -34965, -35581, -27774, -28885, -34788, -26570, -28678, -35188, -35054, -34053, -25933, -34034, -31932, -31466, -32694, -23114, -24503, -23487, -23856, -24795, -26361, -21551, -27304, -26090, -26746, -14429, -13392, -22599, -17422, -14073, -17394, -10667, -11880, -12269, -12998, -5901, -2906, -3684, -6273, 1440, -5475, -795, 5629, -1305, -162, 9368, 372, 4519, 9405, 6082, 12652, 15958, 13719, 16844, 19908, 14424, 20138, 15514, 21621, 26728, 28927, 25005, 23492, 29131, 33411, 29554, 36177, 27797, 27711, 30870, 32940, 34070, 33546, 38909, 32360, 36765, 36095, 36804, 34907, 41272, 37951, 36794, 35261, 38953, 42405, 46445, 36581, 47058, 37754, 46202, 45724, 47011, 37419, 41620, 40136, 37015, 41477, 41422, 36220, 39378, 44463, 37824, 39631, 35504, 30210, 32527, 37824, 31463, 27375, 31581, 28853, 32323, 28678, 30964, 29995, 21282, 19316, 26525, 23094, 14352, 23696, 17824, 16876, 16309, 16839, 16645, 9601, 4651, 11120, 4912, 9671, 2665, 6809, -2405, -4322, 3385, -8024, -1593, -2331, -7196, -9158, -3177, -11409, -12119, -16719, -15834, -17106, -11205, -20080, -20346, -20162, -17519, -25252, -17366, -27719, -23963, -29930, -21938, -23259, -29747, -24724, -26744, -23700, -27669, -23927, -30089, -31127, -29796, -32803, -24830, -30500, -33109, -30963, -27632, -31140, -33637, -25291, -28308, -30533, -32001, -31620, -27502, -28062, -23793, -31278, -21261, -22586, -28398, -18915, -26034, -20257, -20131, -23782, -24695, -14449, -13484, -16551, -19835, -12320, -16118, -8242, -9370, -11523, -2259, -2897, -49, -8606, -5900, 2109, 2967, 5287, 3327, 3767, 7370, 11682, 10813, 10396, 9037, 15267, 12714, 16281, 21451, 22204, 24154, 25897, 25645, 17044, 18255, 20438, 23664, 21904, 27820, 27864, 31291, 36907, 30278, 31657, 38807, 33371, 31712, 36907, 41808, 36762, 41120, 40860, 39229, 39971, 46125, 36045, 38726, 41006, 42914, 46574, 41759, 41437, 45169, 41771, 46414, 41514, 41699, 41323, 37915, 35832, 35216, 44670, 36276, 43312, 40916, 42224, 42331, 31981, 34280, 40546, 35648, 37793, 31871, 25262, 31603, 25845, 28351, 29635, 27090, 25704, 22653, 19164, 20162, 13861, 19808, 22730, 11025, 8984, 17911, 8861, 4641, 13004, 3512, 11064, 241, 1980, 3525, 2072, 1720, 145, -3771, -8625, -2543, -9977, -6314, -5064, -15608, -6103, -18618, -10071, -11186, -21749, -16824, -13057, -21541, -16645, -20033, -18639, -19359, -29193, -27128, -23372, -26012, -20805, -24083, -26787, -30507, -31453, -24232, -29865, -25694, -34578, -25578, -35738, -25306, -25323, -29829, -34622, -33799, -27249, -25509, -34833, -25784, -23001, -29978, -25938, -28972, -29925, -22436, -22533, -27181, -22768, -23920, -27050, -26995, -20448, -22062, -20333, -19942, -20290, -16448, -11732, -16542, -9789, -11282, -10178, -12045, -10563, -4177, -7067, -2248, 3723, 2284, 3206, 7938, 7078, 6419, 11886, 2537, 6418, 16431, 15195, 12956, 16766, 14901, 15762, 15039, 18356, 15347, 21915, 21447, 30376, 26463, 31098, 26912, 28629, 34056, 37044, 32374, 38143, 36784, 35564, 41212, 40239, 42591, 39493, 36911, 38669, 44460, 34137, 36293, 40487, 41695, 36165, 43627, 46616, 37356, 41407, 39550, 48043, 43443, 39051, 37428, 42188, 45334, 45130, 44722, 36717, 40363, 43839, 34190, 42454, 42328, 33411, 30974, 34984, 38512, 33241, 31668, 31801, 26276, 25347, 33203, 28899, 23720, 29811, 18919, 22547, 24521, 18663, 18155, 18394, 21528, 18821, 8949, 10140, 10009, 14509, 7789, 4256, 7207, 4417, 8110, 7188, 4428, 1770, 849, 1413, -9959, -7989, -13264, -4590, -9694, -12612, -15485, -12934, -17030, -20804, -21682, -22927, -19821, -24252, -21337, -16741, -24179, -27816, -23184, -20233, -27275, -31622, -31015, -32365, -24869, -28756, -26616, -26606, -28462, -28035, -25245, -28005, -25547, -30525, -34467, -35307, -27422, -32175, -27600, -27579, -28745, -26178, -28317, -28074, -27461, -21636, -27640, -30287, -28121, -22038, -19411, -17024, -25278, -17816, -19013, -20234, -17942, -17082, -14137, -11926, -16124, -17529, -7468, -11522, -5641, -11575, -11149, -264, 693, 3500, 3197, -5439, 2034, 8851, 4344, 10078, 1756, 14179, 14757, 11788, 11534, 11743, 17687, 10475, 16120, 24019, 20747, 21116, 22612, 21550, 30463, 31985, 27455, 34319, 28903, 29567, 27989, 28700, 37326, 36922, 35384, 39788, 36715, 37907, 34488, 39623, 34830, 34264, 42351, 41880, 37571, 40152, 43129, 42460, 37481, 38112, 36161, 41216, 42039, 37999, 43984, 35980, 36977, 46734, 46689, 34914, 40067, 44037, 36037, 42595, 41727, 38836, 30570, 34369, 39901, 36364, 31852, 33990, 28351, 31320, 35245, 32596, 24680, 28374, 23316, 29724, 17638, 18420, 23941, 13911, 18016, 19964, 17905, 9377, 11611, 9209, 9400, 9354, 2667, 10462, 5902, -1213, 2290, 5350, 2218, -287, -4252, -8040, -5603, -10739, -11140, -5237, -6753, -9028, -8602, -18737, -15751, -15498, -13081, -17086, -21364, -18061, -18014, -21483, -28506, -19175, -30374, -25345, -30901, -28339, -23663, -31015, -23739, -26207, -30588, -32444, -32644, -26638, -35433, -27865, -28692, -27159, -24319, -31362, -32692, -25035, -25632, -29478, -33577, -27457, -31539, -26878, -28450, -28332, -22715, -24565, -20513, -26800, -20267, -26948, -17018, -17557, -13356, -22647, -11752, -15480, -13106, -15572, -17284, -6771, -14070, -10107, -5812, -11, -4507, 2508, -5381, -1979, 2965, -3303, 6290, 3706, 9783, 5941, 6572, 15972, 14094, 11761, 9302, 18293, 18430, 12930, 14770, 26411, 21803, 17298, 18867, 21082, 31294, 27246, 29469, 29714, 25580, 36563, 30159, 30825, 35608, 35004, 34487, 38689, 42791, 39609, 36142, 35763, 39094, 34589, 45239, 42394, 37807, 41885, 36478, 46388, 41444, 42771, 43007, 44333, 40512, 36832, 41195, 36022, 44050, 35259, 45910, 42910, 44768, 39113, 35239, 34834, 40172, 42275, 33832, 37800, 29200, 34183, 31249, 33903, 27242, 24202, 27429, 28611, 21358, 24070, 25291, 26192, 18705, 18590, 23129, 19626, 12790, 17717, 10732, 9229, 4607, 7696, 7086, 4124, 2598, 653, 7664, 5388, -1542, -1888, -2183, -4406, -8356, -959, -11943, -5012, -16231, -13821, -9969, -12375, -19222, -10869, -16856, -21398, -18441, -15331, -16485, -22342, -23657, -26031, -29876, -22162, -30325, -28244, -28335, -22956, -33856, -24363, -31448, -32234, -29645, -26973, -33500, -33464, -24376, -29021, -32478, -24403, -25139, -33472, -35512, -26670, -24459, -33115, -33641, -26421, -25821, -26308, -31826, -22945, -19136, -19257, -27630, -23885, -24367, -19613, -18030, -20802, -13783, -12757, -11844, -15911, -18343, -9278, -4652, -13443, -12788, -1885, -5802, -39, 770, -5417, -3351, -4331, 3712, 7101, 5253, 789, 13760, 9218, 8537, 7980, 14768, 15490, 18929, 13030, 16769, 15474, 25246, 20294, 20745, 18682, 29435, 26891, 28477, 33560, 32809, 33148, 28213, 33622, 39447, 35909, 39280, 42168, 41703, 34278, 32752, 38362, 33630, 39670, 45873, 37802, 39808, 40648, 45711, 45833, 41497, 40717, 47336, 45096, 44997, 47410, 41980, 45164, 40804, 45277, 39382, 43164, 45573, 39599, 37915, 34626, 35378, 32121, 34570, 33244, 32569, 37434, 33090, 32023, 34100, 25202, 30248, 25809, 24555, 26312, 28636, 19422, 23921, 25449, 15718, 15636, 16732, 20166, 14159, 10118, 11873, 11007, 7703, 1541, 8474, 4747, 1872, -3300, -1111, -3954, -5659, 377, -6001, -11393, -8794, -5230, -13819, -6028, -14369, -15407, -18058, -12378, -21863, -12296, -22855, -22285, -18394, -25879, -22269, -20568, -18846, -21956, -22437, -27216, -29844, -27008, -31157, -24103, -26680, -25196, -25779, -29959, -32097, -27701, -24203, -26879, -26168, -27615, -28856, -26811, -29703, -25014, -34328, -23122, -33213, -27362, -28605, -31632, -23602, -24300, -21579, -23465, -19747, -21767, -16490, -16476, -19936, -15581, -18389, -13065, -18103, -9123, -16411, -17731, -8369, -6197, -3868, -9795, -2772, -4688, -4287, 1342, 4254, -4964, 4011, -345, 2992, 2778, 10948, 14274, 11465, 13473, 17573, 15961, 15849, 14903, 19262, 17273, 19073, 19848, 22273, 23894, 29977, 22634, 25346, 29273, 29278, 27592, 32407, 36961, 28019, 33476, 30012, 36582, 37046, 40513, 34727, 39618, 38642, 44016, 42080, 38809, 39108, 38312, 47019, 39359, 37853, 40428, 45091, 44686, 44600, 36147, 40457, 46634, 39372, 42452, 38513, 36049, 38795, 43494, 44939, 42929, 32927, 35324, 33390, 33623, 40867, 34771, 36319, 36521, 27430, 35319, 24674, 31335, 30058, 28796, 20607, 23199, 22760, 21799, 24524, 21065, 21327, 16716, 20522, 8473, 12861, 8381, 9429, 10530, 3420, 6879, 2116, 7443, -2925, -4648, 4341, -6711, -8035, -9303, -11387, -8259, -6924, -6196, -7898, -10016, -14067, -12349, -10439, -16960, -20414, -15569, -23206, -24159, -22269, -21253, -22111, -28818, -29528, -28270, -23463, -27963, -23468, -22682, -29592, -34171, -28261, -26430, -31831, -29945, -33362, -24803, -30356, -29651, -33437, -34835, -35104, -25734, -26049, -32678, -23880, -26009, -25878, -21347, -32325, -27012, -25570, -23748, -29042, -21305, -27813, -20866, -18093, -19856, -17316, -21174, -14921, -17039, -19270, -14831, -15049, -14118, -8301, -8269, -8334, -9413, -393, 946, -4689, 642, 3965, 7431, 8364, 3277, 1961, 10971, 4097, 5998, 9725, 17001, 15140, 16504, 21909, 18974, 13437, 24334, 23153, 22814, 21455, 22495, 26321, 24370, 23292, 25792, 27879, 28126, 33982, 37513, 38218, 38939, 38585, 41147, 40897, 34585, 44709, 34418, 41644, 36855, 37614, 39134, 37738, 41727, 47293, 40750, 43150, 43476, 44789, 40970, 46389, 46988, 44746, 38889, 44756, 36522, 40488, 41322, 41950, 37545, 41121, 42399, 31694, 31964, 39937, 33807, 32832, 38549, 35103, 36921, 26908, 24219, 26629, 26926, 26642, 30386, 23370, 21054, 26987, 16885, 20490, 22806, 17967, 12163, 13629, 5901, 15191, 8054, 5450, 11917, 4645, 1197, -2610, 2036, -4486, -6788, -1996, -6850, -7246, -4153, -3808, -11207, -5028, -6326, -16513, -10881, -13841, -11270, -16141, -15963, -16451, -21726, -24252, -27717, -23303, -22012, -27179, -25007, -28954, -28948, -25265, -22885, -23729, -32010, -30110, -24547, -32440, -24106, -28477, -34078, -26186, -28268, -29559, -33041, -35459, -32950, -31179, -27615, -23031, -32044, -24983, -22947, -27414, -30619, -22138, -25506, -29141, -19231, -21337, -26987, -16330, -25948, -24939, -12509, -15133, -17808, -15181, -10938, -18408, -9071, -8168, -9869, -7136, -8804, -9552, -5497, 2095, -4944, -1978, -1071, -2623, 3910, 9134, 11362, 10543, 7796, 8127, 14224, 17841, 19703, 10854, 16999, 14014, 16788, 25649, 18587, 18890, 25165, 23559, 25500, 31536, 33177, 32295, 30120, 33809, 29565, 35316, 36863, 36778, 34473, 35414, 33767, 41925, 38863, 37740, 43304, 37259, 44988, 44994, 45649, 40156, 40510, 46420, 41722, 43051, 44547, 47690, 42579, 43505, 42500, 46531, 45453, 36722, 36415, 36735, 42354, 35133, 43980, 40035, 32899, 40396, 40231, 40039, 34461, 33466, 27869, 30957, 30365, 24699, 27584, 26973, 21780, 25732, 17345, 19656, 21002, 17257, 19301, 15109, 11063, 19132, 14502, 13378, 12226, 11703, 11518, 6230, 468, 1865, 5817, -3368, -2800, 3541, 287, -8066, 16, -12548, -9444, -10937, -12201, -16869, -14267, -13122, -9715, -20055, -19482, -21553, -22224, -24407, -27305, -23024, -26328, -19571, -24410, -20456, -20384, -25672, -31854, -22626, -27103, -24019, -29919, -28030, -34763, -24678, -28249, -34843, -27719, -31399, -35105, -33448, -32889, -32960, -26969, -26054, -28201, -27730, -26354, -21581, -25274, -25094, -20737, -24137, -26252, -17989, -23417, -20619, -18299, -17872, -22527, -23108, -19749, -11531, -14148, -14163, -13421, -8094, -8335, -7059, -11797, -7254, -5088, -5348, -2763, -3095, 3488, 96, 5402, 3982, 8338, 12214, 8508, 14520, 7615, 16861, 8666, 14608, 10575, 21356, 15054, 16152, 17592, 24962, 20402, 22592, 29409, 27306, 33317, 24104, 29696, 32318, 33184, 37218, 29681, 32615, 29816, 42011, 40492, 40975, 34210, 37320, 35459, 40101, 44292, 42553, 43554, 43245, 44558, 46311, 43631, 38326, 43087, 38121, 46997, 36876, 39846, 42535, 40983, 44633, 40942, 36853, 42189, 34900, 40471, 39561, 34017, 32740, 31797, 30800, 30605, 38799, 26562, 36964, 24739, 35116, 25939, 27594, 30543, 29807, 20103, 24592, 26752, 25923, 14194, 13767, 19312, 9593, 8529, 12229, 15233, 15653, 2324, 7452, 9932, 9145, 7015, 6064, 3114, -5808, -2417, -7838, -1157, -1277, -11695, -4334, -11543, -12814, -15336, -9300, -11952, -16591, -14501, -12706, -22993, -23107, -19255, -18122, -18432, -24730, -28904, -30052, -27353, -22339, -30335, -23926, -26064, -34088, -25326, -24024, -29509, -25636, -34305, -26873, -24966, -26131, -33035, -33534, -29693, -31038, -29839, -23367, -27749, -23280, -28347, -28518, -23972, -23759, -26787, -30839, -29725, -20424, -21361, -28053, -20864, -18000, -24408, -22151, -13972, -21034, -10995, -9384, -19229, -13670, -15004, -9298, -13349, -12843, -787, 970, -5084, -345, -5959, -2927, -3605, 2935, 446, 11953, 24280, 20903, -2456, 57, 23924, 32985, 4998, 2129, 20949, 30619, 33232, 11129, 15115, 29677, 47673, 25995, 4847, 21442, 49328, 45107, 14615, 17072, 36881, 57336, 33128, 22620, 27259, 57337, 46779, 31254, 17305, 46042, 59147, 41479, 20399, 36190, 51306, 55664, 27433, 21151, 44281, 64330, 42327, 28498, 33591, 48490, 56612, 40203, 18390, 43365, 59424, 47287, 23663, 26800, 47474, 48305, 29303, 18248, 34092, 56298, 47487, 13249, 19135, 40074, 45974, 24020, 8576, 23359, 46547, 29133, 13458, 6842, 31396, 31453, 14715, -7271, 7976, 31761, 21677, -3380, -9193, 11781, 27397, 7506, -14861, -1426, 20591, 15181, -14791, -18743, -3425, 18393, -4936, -22008, -19580, -1914, 5761, -25048, -35687, -20712, 6088, -6622, -38276, -32850, -14289, -4020, -21211, -43956, -20122, -9123, -20024, -37824, -34735, -16886, -15666, -31875, -50588, -36631, -18258, -14029, -38580, -46717, -19380, -9292, -28676, -49163, -38398, -19600, -19262, -39549, -46065, -22641, -10298, -22025, -49664, -36230, -11487, -15723, -32594, -47118, -20582, -788, -17636, -38356, -35204, -12695, -34, -20466, -36578, -19874, 2145, -2345, -22945, -20985, 6807, 13580, -16032, -21844, -6780, 9008, 11870, -14272, -9620, 5811, 18095, 4675, -15986, 5019, 24185, 24398, 1375, -3447, 18831, 31742, 22259, 202, 12416, 35738, 40000, 9438, 12884, 24503, 43066, 33495, 9990, 22841, 44491, 40116, 25494, 17925, 38820, 51714, 40743, 23117, 31774, 45379, 49380, 34641, 25404, 46317, 54079, 46201, 28328, 27842, 56932, 55921, 33240, 26231, 36339, 63777, 53763, 26950, 21682, 45868, 55542, 42927, 23459, 33173, 53082, 48612, 30644, 27362, 43535, 55380, 37939, 10965, 27855, 42512, 43216, 19772, 7659, 27989, 50821, 29228, 6604, 13893, 32789, 31553, 10091, 166, 23760, 34666, 19538, -6670, 6835, 25950, 29424, 3983, -4539, 11814, 19420, 11465, -10573, -11809, 14100, 10555, -12437, -28763, -12462, 10326, 296, -25104, -27219, -9462, 7649, -15089, -34274, -24261, 2302, -4196, -27845, -36316, -9218, -533, -28318, -44948, -27584, -11313, -14123, -31889, -38018, -20073, -9281, -21363, -46266, -42064, -17749, -18318, -37973, -52491, -33064, -16109, -20206, -42620, -37954, -11612, -8135, -29900, -50758, -22846, -9795, -25912, -44434, -33921, -11003, -14626, -27075, -37897, -28033, -9898, -15097, -38754, -33196, -10328, -1259, -13566, -33874, -20841, -1663, -4153, -25717, -29908, 1389, 5392, -3812, -22720, -12212, 15915, 10360, -13915, -13086, 4669, 28249, 11212, -4708, 4113, 28652, 27900, 7522, 98, 16447, 36072, 27920, -1550, 10805, 34225, 43999, 19938, 14231, 28319, 50254, 35718, 15733, 15196, 44652, 55262, 30101, 16728, 37094, 48863, 50586, 18027, 24767, 50003, 57658, 37614, 20355, 37678, 62629, 54395, 34798, 21866, 48892, 55243, 42749, 26687, 31191, 60590, 52957, 35734, 22589, 40156, 55239, 37378, 27892, 24592, 47854, 46002, 25146, 13479, 39804, 53281, 35619, 13255, 16834, 42242, 39795, 24016, 10358, 24978, 46888, 35777, 5717, 10444, 31421, 34638, 18513, 5405, 15597, 28384, 17866, -612, -4990, 15578, 26108, 819, -10325, -5644, 13598, 9552, -17332, -11637, 8312, 12664, -9138, -25044, -15378, 9069, 1063, -16581, -23978, -3795, 1330, -16225, -29568, -30273, -9578, -5844, -24779, -40221, -23853, -10530, -14548, -40117, -37779, -11935, -8099, -36101, -43373, -31946, -5474, -19906, -48704, -42735, -17625, -8455, -34244, -46669, -30220, -7769, -25435, -44873, -45784, -18271, -7096, -31024, -42595, -34360, -10292, -17412, -33695, -38597, -14137, -10952, -25899, -36954, -31634, -10997, -8094, -24098, -36957, -11338, 758, -17930, -30551, -16960, 32, -1323, -20316, -22551, -5801, 15258, -4781, -15820, -12694, 7351, 16085, -746, -8021, 11865, 30988, 20191, -750, 2711, 24102, 29529, 6471, 587, 20190, 33830, 33419, 2729, 7658, 30165, 38429, 25862, 7392, 29773, 46130, 44301, 13512, 18707, 41190, 55946, 37163, 22869, 35007, 48585, 46831, 31638, 17655, 42997, 55929, 45794, 19092, 36195, 58990, 56185, 30333, 19757, 45976, 54520, 41375, 21232, 30691, 56181, 61040, 34500, 17622, 38188, 59462, 49605, 21138, 25956, 52200, 54562, 32267, 15469, 31419, 54649, 39836, 17698, 15591, 41000, 47107, 27584, 8764, 20072, 40733, 28861, 8795, 11404, 29811, 39024, 20411, 1230, 12065, 31782, 30066, -4755, -8412, 12249, 21618, 1804, -7724, -3585, 10736, 9388, -7884, -21604, -7122, 11395, -6671, -20890, -14817, -4187, 5286, -17474, -34853, -11096, -1039, -16425, -38576, -28178, -7160, -1472, -25135, -37095, -31635, -8452, -19528, -40054, -35850, -21010, -9208, -36063, -50722, -29365, -16537, -14896, -44069, -43122, -28782, -9527, -30151, -42541, -39236, -16131, -22011, -34531, -46403, -29404, -7848, -25734, -46880, -32736, -8518, -14921, -33521, -42498, -25622, -3704, -12358, -42351, -26149, -6399, -4005, -28228, -37132, -15868, 4047, -8063, -23773, -18375, 4081, 7109, -10106, -21931, -11040, 14189, 4788, -13291, -7543, 10231, 15330, 8031, -6443, 1640, 22679, 24653, -330, -1264, 23471, 28755, 21700, 6070, 8245, 40461, 39567, 6932, 8558, 32105, 43589, 32088, 15055, 22321, 46648, 43348, 28397, 15818, 38605, 57632, 38053, 19488, 27752, 50068, 49284, 35781, 16585, 39586, 53017, 53573, 26472, 34280, 51142, 63065, 34705, 29081, 44683, 58110, 52242, 28737, 32466, 46648, 52286, 43025, 19044, 32253, 57383, 47035, 29702, 26862, 48842, 52525, 38928, 12571, 28461, 50379, 39156, 20537, 18100, 30384, 42511, 32912, 8157, 11342, 33746, 37682, 12649, -366, 21810, 37429, 17319, -3282, 515, 27238, 20988, 6944, -12911, 6024, 25852, 12097, -17548, -9416, 5409, 19659, -3245, -22587, -6114, 15663, -4348, -20678, -20991, -82, 120, -17619, -39506, -23282, -5762, -8699, -31220, -32400, -15861, -4255, -18103, -36972, -30873, -5341, -19121, -33613, -45616, -26543, -6293, -28208, -50244, -43726, -10160, -13690, -34328, -41981, -25694, -7058, -28535, -41721, -35426, -19693, -19289, -32553, -51543, -25616, -10791, -18953, -46150, -38307, -13426, -14485, -29123, -36894, -29614, -5335, -10317, -36439, -27569, -7007, -3363, -17569, -28342, -17537, 6828, 3995, -18450, -28683, -4799, 7152, -10830, -27531, -8021, 15391, 17579, -6320, -15912, 8656, 20710, 12013, -13523, 3913, 28685, 29254, 3021, -1160, 18232, 30714, 27384, 6063, 7994, 40697, 35311, 15956, 7336, 24114, 42469, 38571, 11335, 19335, 40572, 49230, 34819, 13548, 27536, 58677, 48165, 24189, 24894, 43063, 62856, 36174, 24029, 35167, 51711, 52740, 29521, 23647, 43277, 64065, 36756, 22196, 38860, 62940, 55217, 34284, 27662, 47270, 60607, 47699, 22884, 29199, 54556, 51165, 24140, 18637, 38661, 51812, 37461, 19979, 22037, 43713, 40770, 19773, 9981, 28955, 46466, 37625, 13793, 5356, 37531, 32486, 20097, 757, 10940, 27046, 20001, 2205, -8027, 16618, 21065, 549, -17757, 2147, 14231, 13535, -16169, -14641, 4116, 11324, -1163, -20366, -9084, 286, 3883, -27970, -33692, -13980, 1585, -16835, -36086, -29796, -6489, -7043, -27979, -35578, -23199, -1302, -16870, -37425, -40134, -19164, -10291, -31663, -50379, -33248, -9825, -18696, -40895, -46996, -16440, -8770, -35174, -53370, -35520, -10076, -26790, -44647, -43038, -15137, -15317, -35538, -44520, -36989, -5064, -19106, -37198, -36902, -14117, -6383, -20093, -35176, -23375, -8824, -6761, -25932, -37773, -9202, 2157, -11221, -33443, -25909, 504, 9183, -17615, -27269, -573, 16617, -4681, -13868, -7785, 10856, 19256, -5810, -7917, 3400, 21167, 18368, -5436, 932, 29065, 28253, 5859, 2237, 14178, 37574, 25499, 2803, 4944, 36902, 40214, 22883, 11424, 28064, 49357, 39906, 15647, 19203, 34283, 49621, 36966, 19419, 28048, 58675, 45995, 30973, 18811, 43538, 62347, 41281, 18755, 33354, 52855, 51358, 35715, 24760, 40633, 55443, 43057, 21293, 29162, 59536, 57133, 31476, 22307, 42472, 58329, 47466, 28059, 24543, 51362, 49276, 26500, 15575, 36309, 49627, 47425, 19419, 15234, 43996, 51093, 29982, 5938, 18710, 44380, 36516, 9777, 11386, 26138, 42231, 17094, -1822, 11167, 27175, 23730, -4496, -4042, 13131, 26327, 10981, -16815, -2000, 19861, 11126, -7630, -22105, -4755, 8495, -388, -24062, -16036, -1020, -428, -20457, -32176, -11794, -3008, -16129, -32135, -37449, -14096, -2544, -26440, -40505, -22309, -3771, -16487, -42517, -45029, -13704, -4732, -25014, -44898, -38328, -17986, -22702, -47763, -42473, -27675, -10714, -26650, -47087, -38179, -10765, -19706, -42314, -42153, -24350, -13343, -23013, -48871, -30715, -15919, -16972, -39077, -38465, -17664, -2017, -14519, -32060, -31377, -3547, -4063, -18685, -40101, -9430, 4498, -8162, -26373, -25392, -2853, 10230, -9141, -20106, -8374, 11221, 5204, -16305, -7737, 14200, 18406, 4133, -8360, 7522, 30420, 22348, -5672, -5418, 25697, 32635, 19151, 4148, 10069, 36946, 31370, 6879, 11488, 24527, 43685, 27303, 8319, 23365, 50059, 40076, 27271, 20313, 41935, 59333, 36240, 20912, 30980, 52397, 59696, 38224, 27847, 35216, 57843, 45675, 21790, 24934, 56239, 58728, 43016, 30037, 38838, 57781, 47441, 27271, 24890, 49601, 57460, 35537, 17821, 34356, 55766, 47273, 28002, 21550, 42696, 57375, 39100, 19746, 30439, 47995, 44815, 21737, 8567, 30167, 47105, 26465, 11429, 12727, 31440, 33325, 12570, 7800, 22616, 37453, 20675, -1822, 6707, 22556, 24877, -1422, -7272, 6592, 20713, 12386, -18037, -17736, 11055, 16201, -6940, -17824, -6637, 10223, -2731, -29132, -22138, -7524, 1200, -19659, -33083, -20678, 2117, -3646, -28625, -30261, -18746, 545, -28721, -44911, -37336, -8109, -8836, -36461, -47780, -23243, -9363, -30137, -48330, -35431, -15012, -20177, -40119, -48523, -26941, -17886, -24666, -41160, -45232, -14483, -8471, -34464, -43890, -30753, -10656, -26227, -43547, -40354, -17601, -4807, -29363, -37855, -21461, -7259, -17447, -39331, -31341, -10263, 5063, -19226, -37087, -17752, 9056, 1174, -23843, -27138, 3144, 16695, -6633, -26829, -13024, 14990, 8740, -11651, -13977, 6864, 21433, 8722, -12086, -4748, 26861, 22183, 8634, -3279, 16525, 38657, 26391, -111, 6188, 31105, 40661, 22491, 8528, 23261, 48730, 41002, 11793, 23538, 39556, 53739, 34024, 17256, 33280, 58475, 40750, 24123, 26085, 50667, 53609, 32109, 18166, 39703, 63312, 50829, 35361, 24607, 44384, 58555, 42959, 26025, 35944, 55013, 50066, 26742, 20538, 47979, 58198, 37745, 24883, 26565, 56162, 52050, 29151, 15847, 41518, 53396, 39544, 16008, 24434, 38681, 46874, 27142, 9996, 29132, 41571, 32981, 5916, 13885, 35634, 42028, 13753, -932, 15276, 36358, 16759, -5347, 2426, 23774, 24935, 8419, -7305, 1796, 17677, 10989, -12973, -14313, 3711, 19387, -6901, -26146, -9594, 6859, 5196, -26553, -29510, -14366, 5157, -11240, -29179, -24847, -2835, -1826, -30055, -39546, -16735, -1534, -23503, -47077, -41646, -18229, -15584, -32576, -51369, -28708, -8853, -27106, -47870, -44588, -23175, -15765, -30967, -50610, -29077, -12236, -20590, -40955, -40224, -15776, -16170, -27366, -50028, -37947, -15387, -20487, -42962, -35472, -20831, -913, -21571, -35689, -29813, -8559, -11099, -28815, -37041, -14521, -3390, -11170, -24978, -16684, -2995, 5769, -18956, -29143, -3251, 12327, 1298, -13794, -15608, 12189, 11901, -4789, -10420, 1147, 27175, 12957, -3971, -5116, 22672, 24631, 7699, -4127, 15939, 33112, 27462, 10893, 8078, 27604, 41288, 23975, 13529, 21870, 50026, 42215, 14014, 14543, 41343, 51995, 31661, 15161, 33533, 54193, 46247, 30735, 21764, 43872, 60840, 41779, 18009, 27538, 56679, 55143, 38451, 20045, 42957, 60806, 41973, 30575, 32894, 58992, 58320, 28661, 20850, 35753, 59315, 40854, 25778, 25710, 46015, 53612, 34324, 21290, 30263, 48828, 39857, 20155, 21539, 41992, 50821, 30230, 4925, 25519, 46546, 37346, 14389, 531, 28196, 34142, 18900, 2715, 6402, 31741, 20292, 169, -5622, 14924, 22201, 4537, -8428, -4928, 10075, 15174, -14067, -16829, 2381, 10464, -6762, -21293, -22192, -1200, -140, -24824, -31256, -16393, 4461, -10874, -35061, -37059, -13162, -4361, -27707, -36184, -31379, -7993, -16053, -44236, -39949, -14056, -14044, -34503, -51853, -31449, -18663, -21392, -36403, -41994, -26475, -10157, -34512, -46321, -32396, -9822, -19182, -40301, -43425, -21933, -10933, -27453, -47456, -40903, -13238, -15982, -35157, -36644, -21358, 78, -22554, -31676, -35838, -9260, 312, -22801, -34499, -17668, -772, -8782, -31086, -25183, -3446, 12241, -5675, -27029, -4063, 8676, 8476, -12196, -18472, 5123, 16648, 7223, -14268, 3731, 25841, 22010, -2482, -3062, 20210, 39505, 11875, -518, 16622, 37426, 32334, 17670, 3367, 28110, 49640, 32186, 14110, 21094, 40732, 51459, 28913, 15946, 41057, 51502, 39228, 24239, 22266, 56192, 48212, 30368, 16776, 39742, 62091, 52822, 26604, 33007, 53305, 61454, 31742, 23869, 36914, 57018, 56365, 24411, 27955, 46785, 59079, 44443, 17799, 40812, 51148, 45608, 27542, 17752, 38423, 55762, 29596, 22556, 27426, 46458, 46643, 25556, 11995, 35559, 46940, 32136, 9318, 14041, 41221, 32471, 15471, 8135, 17698, 37363, 21948, -3251, 2155, 29260, 30847, 4904, -11765, 483, 23432, 10743, -15071, -7202, 11384, 15777, -10368, -27896, -10765, 6716, -1690, -19518, -29030, -7601, 3952, -15513, -37734, -19542, 2791, -4699, -34931, -38156, -18713, -5281, -25326, -44439, -26207, -11387, -15171, -36214, -48828, -26826, -7484, -25472, -49825, -33895, -16570, -15324, -38339, -51073, -32911, -12524, -31262, -47155, -39794, -15609, -19761, -33246, -50526, -27249, -8859, -17492, -47515, -34409, -16435, -9836, -30871, -40885, -27427, -6256, -14061, -32394, -31017, -3416, 5531, -20034, -36617, -13175, 1237, -153, -17516, -29175, -3973, 10449, -4212, -16794, -12582, 19708, 11731, -5702, -13210, 6675, 22801, 11832, -3883, 5649, 20545, 21714, 9729, -331, 13063, 35747, 28176, 2443, 8292, 31828, 35519, 16925, 9550, 24499, 47623, 39767, 10412, 21830, 44822, 49374, 34911, 12108, 34748, 50561, 40355, 24972, 28754, 48537, 60963, 34316, 23981, 32522, 55110, 46388, 31841, 32152, 51761, 63040, 42711, 21783, 32366, 54667, 59759, 27684, 25366, 41892, 57827, 38094, 20961, 33963, 56273, 56751, 29054, 23203, 40600, 47569, 34418, 13732, 18713, 39853, 42535, 20070, 16058, 25443, 41496, 30533, 6197, 13375, 30371, 32029, 15837, -2155, 12420, 27024, 26839, -2084, -8016, 23256, 22870, 6044, -10525, -3904, 24763, 14117, -11738, -12018, 4820, 8151, -5358, -20491, -11522, 7183, -3730, -19397, -29556, -7314, 6240, -10021, -39909, -23403, -4315, -11202, -32663, -43465, -19649, -4956, -24968, -35468, -39303, -16149, -14026, -39615, -45359, -31317, -12106, -17065, -39632, -46612, -18120, -15332, -31953, -47910, -35284, -12955, -16958, -41031, -47151, -24742, -13369, -26543, -44055, -30650, -15219, -21144, -33945, -41680, -18245, -6729, -23047, -42930, -31447, -561, -2401, -28116, -35713, -10990, 4483, -7467, -35532, -20432, 2075, 5566, -16549, -27795, -8512, 7426, -4224, -20588, -8011, 10992, 18660, 2589, -11316, 6509);
end;
