-- W2000 definitions
  constant  CFG_DSO_ENABLE             : integer := CONFIG_DSO_ENABLE;
  constant  CFG_DSO_PLATTFORM          : integer := CONFIG_DSO_PLATTFORM;
  constant  CFG_DSO_CHANNELS           : integer := CONFIG_DSO_CHANNELS;
  constant  CFG_DSO_SAMPLING_FREQUENCY : integer := CONFIG_DSO_SAMPLING_FREQUENCY;
  constant  CFG_DSO_INPUT_BIT_WIDTH    : integer := CONFIG_DSO_INPUT_BIT_WIDTH;

