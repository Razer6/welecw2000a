------------------------------------------------------------------------
-- Script created table file
------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library DSO;
use DSO.Global.all;

package pFirCoeff is
constant cFirCoeff : aInputValues(0 to 128-1) := ( 118, -44, -1500, 6464, 11102, 1072, -1142, 314, 314, -1142, 1072, 11102, 6464, -1500, -44, 118, 56, 78, -861, 2530, 5799, 1146, -760, 191, 130, -159, -623, 3957, 5133, 49, -475, 193, 193, -475, 49, 5133, 3957, -623, -159, 130, 191, -760, 1146, 5799, 2530, -861, 78, 56, -111, 22, 1828, 1656, -75, 0, 0, 0, -144, 144, 1974, 1465, -147, 0, 0, 0, -176, 290, 2089, 1261, -195, 0, 0, 0, -203, 458, 2169, 1052, -221, 0, 0, 0, -222, 644, 2209, 844, -229, 0, 0, 0, -229, 844, 2209, 644, -222, 0, 0, 0, -221, 1052, 2169, 458, -203, 0, 0, 0, -195, 1261, 2089, 290, -176, 0, 0, 0, -147, 1465, 1974, 144, -144, 0, 0, 0, -75, 1656, 1828, 22, -111, 0, 0, 0);
end;
