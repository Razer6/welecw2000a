
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
  generic (
    gAddrWidth : integer := 14);
  port (
    iClk  : in  std_ulogic;
    oData : out std_ulogic_vector(31 downto 0);
    iAddr : in  std_ulogic_vector(31 downto 0));
end entity;

architecture Rtl of ROM is
  subtype aDataVec is std_ulogic_vector(31 downto 0);
  type    aMem is array (2**gAddrWidth-1 downto 0) of aDataVec;

  constant mem : aMem := (
     0 => x"7f454c46",
     1 => x"01020100",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"0002006a",
     5 => x"00000001",
     6 => x"00000000",
     7 => x"00000034",
     8 => x"00000134",
     9 => x"00000000",
    10 => x"00340020",
    11 => x"00020028",
    12 => x"000b0008",
    13 => x"00000001",
    14 => x"00000074",
    15 => x"00000000",
    16 => x"00000000",
    17 => x"00000065",
    18 => x"00000065",
    19 => x"00000005",
    20 => x"00000001",
    21 => x"00000001",
    22 => x"000000d9",
    23 => x"00000068",
    24 => x"00000068",
    25 => x"00000008",
    26 => x"00000008",
    27 => x"00000006",
    28 => x"00000001",
    29 => x"0b0b0b0b",
    30 => x"80700b0b",
    31 => x"0b80ec0c",
    32 => x"3a0b0b0b",
    33 => x"80de0400",
    34 => x"00000000",
    35 => x"00000000",
    36 => x"00000000",
    37 => x"803d0d80",
    38 => x"51830b86",
    39 => x"8da00c70",
    40 => x"802e8838",
    41 => x"70812e8d",
    42 => x"38963981",
    43 => x"0b868da0",
    44 => x"0c8151eb",
    45 => x"3981c70b",
    46 => x"868da00c",
    47 => x"8251e039",
    48 => x"800b868d",
    49 => x"a00c8111",
    50 => x"51847125",
    51 => x"d238823d",
    52 => x"0d04c13f",
    53 => x"800b800c",
    54 => x"04000000",
    55 => x"00000000",
    56 => x"00002e73",
    57 => x"796d7461",
    58 => x"62002e73",
    59 => x"74727461",
    60 => x"62002e73",
    61 => x"68737472",
    62 => x"74616200",
    63 => x"2e666978",
    64 => x"65645f76",
    65 => x"6563746f",
    66 => x"7273002e",
    67 => x"74657874",
    68 => x"002e6461",
    69 => x"7461002e",
    70 => x"63746f72",
    71 => x"73002e64",
    72 => x"746f7273",
    73 => x"002e6273",
    74 => x"73002e73",
    75 => x"7461636b",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"00000000",
    81 => x"00000000",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"0000001b",
    88 => x"00000001",
    89 => x"00000002",
    90 => x"00000000",
    91 => x"00000074",
    92 => x"00000020",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000020",
    96 => x"00000000",
    97 => x"0000002a",
    98 => x"00000001",
    99 => x"00000006",
   100 => x"00000020",
   101 => x"00000094",
   102 => x"00000045",
   103 => x"00000000",
   104 => x"00000000",
   105 => x"00000001",
   106 => x"00000000",
   107 => x"00000030",
   108 => x"00000001",
   109 => x"00000003",
   110 => x"00000068",
   111 => x"000000d9",
   112 => x"00000008",
   113 => x"00000000",
   114 => x"00000000",
   115 => x"00000001",
   116 => x"00000000",
   117 => x"00000036",
   118 => x"00000001",
   119 => x"00000001",
   120 => x"00000070",
   121 => x"000000e1",
   122 => x"00000000",
   123 => x"00000000",
   124 => x"00000000",
   125 => x"00000001",
   126 => x"00000000",
   127 => x"0000003d",
   128 => x"00000001",
   129 => x"00000001",
   130 => x"00000070",
   131 => x"000000e1",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000001",
   136 => x"00000000",
   137 => x"00000044",
   138 => x"00000008",
   139 => x"00000001",
   140 => x"00000070",
   141 => x"000000e1",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"00000000",
   145 => x"00000001",
   146 => x"00000000",
   147 => x"00000049",
   148 => x"00000001",
   149 => x"00000001",
   150 => x"00ff0000",
   151 => x"000000e1",
   152 => x"00000000",
   153 => x"00000000",
   154 => x"00000000",
   155 => x"00000001",
   156 => x"00000000",
   157 => x"00000011",
   158 => x"00000003",
   159 => x"00000000",
   160 => x"00000000",
   161 => x"000000e1",
   162 => x"00000050",
   163 => x"00000000",
   164 => x"00000000",
   165 => x"00000001",
   166 => x"00000000",
   167 => x"00000001",
   168 => x"00000002",
   169 => x"00000000",
   170 => x"00000000",
   171 => x"000002ec",
   172 => x"00000280",
   173 => x"0000000a",
   174 => x"00000015",
   175 => x"00000004",
   176 => x"00000010",
   177 => x"00000009",
   178 => x"00000003",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"0000056c",
   182 => x"0000010b",
   183 => x"00000000",
   184 => x"00000000",
   185 => x"00000001",
   186 => x"00000000",
   187 => x"00000000",
   188 => x"00000000",
   189 => x"00000000",
   190 => x"00000000",
   191 => x"00000000",
   192 => x"00000000",
   193 => x"00000000",
   194 => x"03000001",
   195 => x"00000000",
   196 => x"00000020",
   197 => x"00000000",
   198 => x"03000002",
   199 => x"00000000",
   200 => x"00000068",
   201 => x"00000000",
   202 => x"03000003",
   203 => x"00000000",
   204 => x"00000070",
   205 => x"00000000",
   206 => x"03000004",
   207 => x"00000000",
   208 => x"00000070",
   209 => x"00000000",
   210 => x"03000005",
   211 => x"00000000",
   212 => x"00000070",
   213 => x"00000000",
   214 => x"03000006",
   215 => x"00000000",
   216 => x"00ff0000",
   217 => x"00000000",
   218 => x"03000007",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"03000008",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"03000009",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"0300000a",
   231 => x"00000001",
   232 => x"00000000",
   233 => x"00000000",
   234 => x"0400fff1",
   235 => x"00000008",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"0400fff1",
   239 => x"00000017",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"0400fff1",
   243 => x"00000022",
   244 => x"00000001",
   245 => x"00000000",
   246 => x"0000fff1",
   247 => x"00000030",
   248 => x"00000000",
   249 => x"00000000",
   250 => x"0400fff1",
   251 => x"00000022",
   252 => x"00000001",
   253 => x"00000000",
   254 => x"0000fff1",
   255 => x"0000003d",
   256 => x"00000037",
   257 => x"00000000",
   258 => x"00000002",
   259 => x"00000041",
   260 => x"00000041",
   261 => x"00000000",
   262 => x"00000002",
   263 => x"00000045",
   264 => x"0000004c",
   265 => x"00000000",
   266 => x"00000002",
   267 => x"00000049",
   268 => x"0000002b",
   269 => x"00000000",
   270 => x"00000002",
   271 => x"0000004e",
   272 => x"00000070",
   273 => x"00000000",
   274 => x"1000fff1",
   275 => x"00000059",
   276 => x"00000070",
   277 => x"00000000",
   278 => x"1000fff1",
   279 => x"00000067",
   280 => x"00000070",
   281 => x"00000000",
   282 => x"1000fff1",
   283 => x"00000073",
   284 => x"00000068",
   285 => x"00000000",
   286 => x"10000003",
   287 => x"0000007d",
   288 => x"00000000",
   289 => x"00000000",
   290 => x"10000001",
   291 => x"00000084",
   292 => x"00000070",
   293 => x"00000000",
   294 => x"10000005",
   295 => x"0000008d",
   296 => x"00000020",
   297 => x"00000056",
   298 => x"12000002",
   299 => x"00000098",
   300 => x"00000070",
   301 => x"00000000",
   302 => x"1000fff1",
   303 => x"000000a4",
   304 => x"00000000",
   305 => x"00000000",
   306 => x"1000fff1",
   307 => x"000000ab",
   308 => x"00000070",
   309 => x"00000000",
   310 => x"1000fff1",
   311 => x"000000b3",
   312 => x"00000070",
   313 => x"00000000",
   314 => x"10000004",
   315 => x"000000c0",
   316 => x"00000070",
   317 => x"00000000",
   318 => x"10000004",
   319 => x"000000c9",
   320 => x"0000005e",
   321 => x"0000000b",
   322 => x"12000002",
   323 => x"000000d2",
   324 => x"00000070",
   325 => x"00000000",
   326 => x"1000fff1",
   327 => x"000000d9",
   328 => x"0000006c",
   329 => x"00000000",
   330 => x"10000003",
   331 => x"000000e5",
   332 => x"00000070",
   333 => x"00000000",
   334 => x"1000fff1",
   335 => x"000000ea",
   336 => x"00ff0000",
   337 => x"00000000",
   338 => x"10000007",
   339 => x"000000f1",
   340 => x"00000068",
   341 => x"00000000",
   342 => x"10000003",
   343 => x"000000fe",
   344 => x"00000070",
   345 => x"00000000",
   346 => x"10000005",
   347 => x"00637274",
   348 => x"302e5300",
   349 => x"3c636f6d",
   350 => x"6d616e64",
   351 => x"206c696e",
   352 => x"653e003c",
   353 => x"6275696c",
   354 => x"742d696e",
   355 => x"3e004f50",
   356 => x"54494d49",
   357 => x"5a455f53",
   358 => x"495a4500",
   359 => x"626f6f74",
   360 => x"6c6f6164",
   361 => x"65722e63",
   362 => x"002e4c36",
   363 => x"002e4c37",
   364 => x"002e4c38",
   365 => x"002e4c31",
   366 => x"35005f62",
   367 => x"73735f65",
   368 => x"6e645f5f",
   369 => x"005f5f62",
   370 => x"73735f73",
   371 => x"74617274",
   372 => x"5f5f005f",
   373 => x"5f627373",
   374 => x"5f656e64",
   375 => x"5f5f005f",
   376 => x"68617264",
   377 => x"77617265",
   378 => x"005f7374",
   379 => x"61727400",
   380 => x"5f5f5f64",
   381 => x"746f7273",
   382 => x"00426f6f",
   383 => x"746c6f61",
   384 => x"64657200",
   385 => x"5f5f6273",
   386 => x"735f7374",
   387 => x"61727400",
   388 => x"5a50555f",
   389 => x"4944005f",
   390 => x"5f656e64",
   391 => x"5f5f005f",
   392 => x"5f5f6374",
   393 => x"6f72735f",
   394 => x"656e6400",
   395 => x"5f5f5f63",
   396 => x"746f7273",
   397 => x"005f7072",
   398 => x"656d6169",
   399 => x"6e005f65",
   400 => x"64617461",
   401 => x"005f6370",
   402 => x"755f636f",
   403 => x"6e666967",
   404 => x"005f656e",
   405 => x"64005f73",
   406 => x"7461636b",
   407 => x"005f5f64",
   408 => x"6174615f",
   409 => x"73746172",
   410 => x"74005f5f",
   411 => x"5f64746f",
   412 => x"72735f65",
   413 => x"6e640065",
others => (others => '-'));
begin  -- Rtl
  wrt : process (iClk)
  begin  -- process write
    if iClk'event and iClk = '0' then   -- FALLING clock edge
      oData <= mem(to_integer(unsigned(iAddr(2**gAddrWidth-1 downto 0))));
    end if;
  end process wrt;
end architecture;
