------------------------------------------------------------------------
-- Script created table file
------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Global.all;

package pFastFirCoeff is
  constant cFastFirCoeff : aInputValues(0 to 128-1) := (
    1, 0, -16, 67, 116, 11, -12, 3,
    3, -12, 11, 116, 67, -16, 0, 1,
    1, 1, -9, 26, 60, 12, -8, 2,
    1, -2, -6, 41, 53, 1, -5, 2,
    2, -5, 1, 53, 41, -6, -2, 1,
    2, -8, 12, 60, 26, -9, 1, 1,
    -1, 0, 19, 17, -1, 0, 0, 0,
    -2, 2, 21, 15, -2, 0, 0, 0,
    -2, 3, 22, 13, -2, 0, 0, 0,
    -2, 5, 23, 11, -2, 0, 0, 0,
    -2, 7, 23, 9, -2, 0, 0, 0,
    -2, 9, 23, 7, -2, 0, 0, 0,
    -2, 11, 23, 5, -2, 0, 0, 0,
    -2, 13, 22, 3, -2, 0, 0, 0,
    -2, 15, 21, 2, -2, 0, 0, 0,
    -1, 17, 19, 0, -1, 0, 0, 0);
end;
