------------------------------------------------------------------------
-- Script created table file
------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library DSO;
use DSO.Global.all;

package pFastFirCoeff is
constant cFastFirCoeff : aInputValues(0 to 128-1) := ( 4, 11, 19, 26, 34, 41, 49, 56, 8, 15, 23, 30, 38, 45, 53, 60, 1, 5, 9, 13, 16, 20, 24, 28, 2, 6, 10, 14, 17, 21, 25, 29, 3, 7, 11, 15, 18, 22, 26, 30, 4, 8, 12, 16, 19, 23, 27, 31, 0, 4, 8, 12, 16, 0, 0, 0, 1, 5, 9, 13, 17, 0, 0, 0, 1, 5, 9, 13, 17, 0, 0, 0, 2, 6, 10, 14, 18, 0, 0, 0, 2, 6, 10, 14, 18, 0, 0, 0, 2, 6, 10, 14, 18, 0, 0, 0, 3, 7, 11, 15, 19, 0, 0, 0, 3, 7, 11, 15, 19, 0, 0, 0, 4, 8, 12, 16, 20, 0, 0, 0, 4, 8, 12, 16, 20, 0, 0, 0);
end;
