------------------------------------------------------------------------
-- Script created table file
------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library DSO;
use DSO.Global.all;

package pFirCoeff is
constant cFirCoeff : aInputValues(0 to 128-1) := ( 964, 2891, 4819, 6746, 8674, 10601, 12529, 14456, 1928, 3855, 5783, 7710, 9638, 11565, 13493, 15420, 248, 1241, 2234, 3227, 4220, 5213, 6206, 7199, 496, 1489, 2482, 3475, 4468, 5461, 6454, 7447, 745, 1738, 2731, 3724, 4717, 5710, 6703, 7696, 993, 1986, 2979, 3972, 4965, 5958, 6951, 7944, 103, 1131, 2159, 3187, 4215, 0, 0, 0, 206, 1234, 2262, 3290, 4318, 0, 0, 0, 308, 1336, 2364, 3392, 4420, 0, 0, 0, 411, 1439, 2467, 3495, 4523, 0, 0, 0, 514, 1542, 2570, 3598, 4626, 0, 0, 0, 617, 1645, 2673, 3701, 4729, 0, 0, 0, 720, 1748, 2776, 3804, 4832, 0, 0, 0, 822, 1850, 2878, 3906, 4934, 0, 0, 0, 925, 1953, 2981, 4009, 5037, 0, 0, 0, 1028, 2056, 3084, 4112, 5140, 0, 0, 0);
end;
